LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY WB_stage IS
    PORT (
        MemtoReg,reset : IN STD_LOGIC;
        ALU_out, MEM_out : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        Result : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END WB_stage;

ARCHITECTURE arch_WB_stage OF WB_stage IS
BEGIN

    Result <= x"00000000" WHEN reset = '1' ELSE ALU_out WHEN MemtoReg = '0' ELSE
        MEM_OUT;

END arch_WB_stage;